module comparator_32 (
    input  wire [31:0] A,  // First 32-bit operand
    input  wire [31:0] B,  // Second 32-bit operand
    output reg is_equal   // Output: 1 if A == B, else 0
);

    // Compute equality using XOR and reduction OR
	 
	 

endmodule